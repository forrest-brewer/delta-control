// --------------------------------------------------------------------
// Copyright 2022 qaztronic
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
//
// Licensed under the Solderpad Hardware License v 2.1 (the "License");
// you may not use this file except in compliance with the License, or,
// at your option, the Apache License version 2.0. You may obtain a copy
// of the License at
//
// https://solderpad.org/licenses/SHL-2.1/
//
// Unless required by applicable law or agreed to in writing, any work
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or
// implied. See the License for the specific language governing
// permissions and limitations under the License.
// --------------------------------------------------------------------

package sd_filter_pkg;

  // --------------------------------------------------------------------
  typedef struct packed {
    int  IN_W ;  // previous node width
    int  IN_N ;  // previous node fractional width
    int  S    ;  // accumulator width
    int  C_W  ;  // accumulator fractional width
    int  C_N  ;  // right shift
    int  OUT_W;  // coefficient width
    int  OUT_N;  // coefficient fractional width
  } sd_filter_cfg_t;

// --------------------------------------------------------------------
endpackage
